
`ifndef APB_SLAVE_SEQUENCER_SV
`define APB_SLAVE_SEQUENCER_SV

function apb_slave_sequencer::new (string name, uvm_component parent);
  super.new(name, parent);
endfunction : new

`endif // APB_SLAVE_SEQUENCER_SV


